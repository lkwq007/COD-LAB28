library verilog;
use verilog.vl_types.all;
entity Decode is
    generic(
        R_type_op       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADD_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ADDU_funct      : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1);
        AND_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        XOR_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        OR_funct        : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        NOR_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        SUB_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0);
        SUBU_funct      : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        SLT_funct       : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi0);
        SLTU_funct      : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        SLL_funct       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SLLV_funct      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        SRL_funct       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        SRLV_funct      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        SRA_funct       : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        SRAV_funct      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        JR_funct        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        BEQ_op          : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        BNE_op          : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        BGEZ_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        BGEZ_rt         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        BGTZ_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        BGTZ_rt         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        BLEZ_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        BLEZ_rt         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        BLTZ_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        BLTZ_rt         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        J_op            : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        ADDI_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        ADDIU_op        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        ANDI_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        XORI_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        ORI_op          : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1);
        SLTI_op         : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        SLTIU_op        : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        SW_op           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1);
        LW_op           : vl_logic_vector(0 to 5) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        alu_add         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        alu_and         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        alu_xor         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        alu_or          : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        alu_nor         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi0);
        alu_sub         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi0, Hi1);
        alu_andi        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi0);
        alu_xori        : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi1, Hi1, Hi1);
        alu_ori         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi0);
        alu_jr          : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi0, Hi1);
        alu_beq         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        alu_bne         : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi0, Hi1, Hi1);
        alu_bgez        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi0);
        alu_bgtz        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi0, Hi1);
        alu_blez        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi0);
        alu_bltz        : vl_logic_vector(0 to 4) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        alu_sll         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi0);
        alu_srl         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi0, Hi1);
        alu_sra         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi0);
        alu_slt         : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi0, Hi1, Hi1);
        alu_sltu        : vl_logic_vector(0 to 4) := (Hi1, Hi0, Hi1, Hi0, Hi0)
    );
    port(
        MemtoReg        : out    vl_logic;
        RegWrite        : out    vl_logic;
        MemWrite        : out    vl_logic;
        MemRead         : out    vl_logic;
        ALUCode         : out    vl_logic_vector(4 downto 0);
        ALUSrcA         : out    vl_logic;
        ALUSrcB         : out    vl_logic;
        RegDst          : out    vl_logic;
        J               : out    vl_logic;
        JR              : out    vl_logic;
        Instruction     : in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of R_type_op : constant is 1;
    attribute mti_svvh_generic_type of ADD_funct : constant is 1;
    attribute mti_svvh_generic_type of ADDU_funct : constant is 1;
    attribute mti_svvh_generic_type of AND_funct : constant is 1;
    attribute mti_svvh_generic_type of XOR_funct : constant is 1;
    attribute mti_svvh_generic_type of OR_funct : constant is 1;
    attribute mti_svvh_generic_type of NOR_funct : constant is 1;
    attribute mti_svvh_generic_type of SUB_funct : constant is 1;
    attribute mti_svvh_generic_type of SUBU_funct : constant is 1;
    attribute mti_svvh_generic_type of SLT_funct : constant is 1;
    attribute mti_svvh_generic_type of SLTU_funct : constant is 1;
    attribute mti_svvh_generic_type of SLL_funct : constant is 1;
    attribute mti_svvh_generic_type of SLLV_funct : constant is 1;
    attribute mti_svvh_generic_type of SRL_funct : constant is 1;
    attribute mti_svvh_generic_type of SRLV_funct : constant is 1;
    attribute mti_svvh_generic_type of SRA_funct : constant is 1;
    attribute mti_svvh_generic_type of SRAV_funct : constant is 1;
    attribute mti_svvh_generic_type of JR_funct : constant is 1;
    attribute mti_svvh_generic_type of BEQ_op : constant is 1;
    attribute mti_svvh_generic_type of BNE_op : constant is 1;
    attribute mti_svvh_generic_type of BGEZ_op : constant is 1;
    attribute mti_svvh_generic_type of BGEZ_rt : constant is 1;
    attribute mti_svvh_generic_type of BGTZ_op : constant is 1;
    attribute mti_svvh_generic_type of BGTZ_rt : constant is 1;
    attribute mti_svvh_generic_type of BLEZ_op : constant is 1;
    attribute mti_svvh_generic_type of BLEZ_rt : constant is 1;
    attribute mti_svvh_generic_type of BLTZ_op : constant is 1;
    attribute mti_svvh_generic_type of BLTZ_rt : constant is 1;
    attribute mti_svvh_generic_type of J_op : constant is 1;
    attribute mti_svvh_generic_type of ADDI_op : constant is 1;
    attribute mti_svvh_generic_type of ADDIU_op : constant is 1;
    attribute mti_svvh_generic_type of ANDI_op : constant is 1;
    attribute mti_svvh_generic_type of XORI_op : constant is 1;
    attribute mti_svvh_generic_type of ORI_op : constant is 1;
    attribute mti_svvh_generic_type of SLTI_op : constant is 1;
    attribute mti_svvh_generic_type of SLTIU_op : constant is 1;
    attribute mti_svvh_generic_type of SW_op : constant is 1;
    attribute mti_svvh_generic_type of LW_op : constant is 1;
    attribute mti_svvh_generic_type of alu_add : constant is 1;
    attribute mti_svvh_generic_type of alu_and : constant is 1;
    attribute mti_svvh_generic_type of alu_xor : constant is 1;
    attribute mti_svvh_generic_type of alu_or : constant is 1;
    attribute mti_svvh_generic_type of alu_nor : constant is 1;
    attribute mti_svvh_generic_type of alu_sub : constant is 1;
    attribute mti_svvh_generic_type of alu_andi : constant is 1;
    attribute mti_svvh_generic_type of alu_xori : constant is 1;
    attribute mti_svvh_generic_type of alu_ori : constant is 1;
    attribute mti_svvh_generic_type of alu_jr : constant is 1;
    attribute mti_svvh_generic_type of alu_beq : constant is 1;
    attribute mti_svvh_generic_type of alu_bne : constant is 1;
    attribute mti_svvh_generic_type of alu_bgez : constant is 1;
    attribute mti_svvh_generic_type of alu_bgtz : constant is 1;
    attribute mti_svvh_generic_type of alu_blez : constant is 1;
    attribute mti_svvh_generic_type of alu_bltz : constant is 1;
    attribute mti_svvh_generic_type of alu_sll : constant is 1;
    attribute mti_svvh_generic_type of alu_srl : constant is 1;
    attribute mti_svvh_generic_type of alu_sra : constant is 1;
    attribute mti_svvh_generic_type of alu_slt : constant is 1;
    attribute mti_svvh_generic_type of alu_sltu : constant is 1;
end Decode;
